/*
   Copyright 2013 Ray Salemi

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/
// vsim -c -do run.do
// vsim -c -do run.do
module top;
   import uvm_pkg::*;
   import   tb_pkg::*;

`include "uvm_macros.svh"


initial begin
   //uvm_config_db #(virtual tinyalu_bfm)::set(null, "*", "bfm", bfm);
   fill_si_array( );
   run_test("test");
end

endmodule : top

     
   