`include "add.svh"
`include "test.svh"
`include "jal.svh"