package OP_pkg;
   import uvm_pkg::*;
`include "uvm_macros.svh"
   `ifdef riscy
      typedef enum bit[31:0] {
                              //no op =32'b00000001000000000000000000000000
                              lsb = 32'b11?????001001?????1?????????????,
                              lsh = 32'b11?????001010?????1?????????????,
                              lub = 32'b11?????000001?????1?????????????,
                              luh = 32'b11?????000010?????1?????????????,
                              lw = 32'b11?????000000?????1?????????????,
                              luw = 32'b00000001000000000000000000000000,
                              LD = 32'b11?????000011?????1?????????????,
                              LSBfAs = 32'b11?????011001?????000001111?????,
                              LSHfAs = 32'b11?????011010?????000001111?????,
                              LUBfAs = 32'b11?????010001?????000001111?????,
                              LUHfAs = 32'b11?????010010?????000001111?????,
                              LWfAs = 32'b11?????010000?????000001111?????,
                              LDfAs = 32'b11?????010011?????000001111?????,
                              LFR = 32'b11?????100000?????1?????????????,
                              LDFR = 32'b11?????100011?????1?????????????,
                              LFSR = 32'b11?????100001?????1?????????????,
                              LCR = 32'b00000001000000000000000000000000,
                              LDCR = 32'b00000001000000000000000000000000,
                              LCSR = 32'b00000001000000000000000000000000,
                              lmorfsm = 32'b00000001000000000000000000000000,
                              lmfps = 32'b00000001000000000000000000000000,
                           lmor&Pfsm = 32'b00000001000000000000000000000000,
                           SB = 32'b11?????001001?????1?????????????,
                           SBiAs = 32'b11?????001001?????1?????????????,
                           SH = 32'b11?????001001?????1?????????????,
                           SHiAs = 32'b11?????001001?????1?????????????,
                           SW = 32'b11?????001001?????1?????????????,
                           SWiAs = 32'b11?????001001?????1?????????????,
                           SD = 32'b11?????001001?????1?????????????,
                           SDiAs = 32'b11?????001001?????1?????????????,
                           SF = 32'b11?????001001?????1?????????????,
                           SDF = 32'b11?????001001?????1?????????????,
                           SFSR = 32'b11?????001001?????1?????????????,
                           SDFdQ = 32'b11?????001001?????1?????????????,
                           SC = 32'b11?????001001?????1?????????????,
                           SDC = 32'b11?????001001?????1?????????????,
                           SCSR = 32'b11?????001001?????1?????????????,
                           SDCdQ = 32'b11?????001001?????1?????????????,
                           Sm = 32'b11?????001001?????1?????????????,
                           SB = 32'b11?????001001?????1?????????????,
                           ALUB = 32'b11?????001001?????1?????????????,
                           ALUBas = 32'b11?????001001?????1?????????????,
                           SRwM = 32'b11?????001001?????1?????????????,
                           Sabbram = 32'b11?????001001?????1?????????????,
                           SRwM(as = 32'b11?????001001?????1?????????????,
                           = 32'b11?????001001?????1?????????????,
                           UIM = 32'b11?????001001?????1?????????????,
                           UIMi = 32'b11?????001001?????1?????????????,
                           UIMami = 32'b11?????001001?????1?????????????,
                           UIMiami = 32'b11?????001001?????1?????????????,
                           SIM = 32'b11?????001001?????1?????????????,
                           SIMi = 32'b11?????001001?????1?????????????,
                           SIMami = 32'b11?????001001?????1?????????????,
                           SIMiami = 32'b11?????001001?????1?????????????,
                           h = 32'b11?????001001?????1?????????????,
                           h( = 32'b11?????001001?????1?????????????,
                           h( = 32'b11?????001001?????1?????????????,
                           A = 32'b11?????001001?????1?????????????,
                           UId = 32'b11?????001001?????1?????????????,
                           UIdi = 32'b11?????001001?????1?????????????,
                           UIdami = 32'b11?????001001?????1?????????????,
                           UIdiami = 32'b11?????001001?????1?????????????,
                           SId = 32'b11?????001001?????1?????????????,
                           SIdi = 32'b11?????001001?????1?????????????,
                           SIdami = 32'b11?????001001?????1?????????????,
                           SIdiami = 32'b11?????001001?????1?????????????,
                           R = 32'b11?????001001?????1?????????????,
                           Ru = 32'b11?????001001?????1?????????????,
                           A = 32'b11?????001001?????1?????????????,
                           Ai = 32'b11?????001001?????1?????????????,
                           Aami = 32'b11?????001001?????1?????????????,
                           Aiami = 32'b11?????001001?????1?????????????,
                           Awc = 32'b11?????001001?????1?????????????,
                           Aiwc = 32'b11?????001001?????1?????????????,
                           Awcami = 32'b11?????001001?????1?????????????,
                           Aiwcami = 32'b11?????001001?????1?????????????,
                           TAami = 32'b11?????001001?????1?????????????,
                           TAiami = 32'b11?????001001?????1?????????????,
                           TAmiatoo = 32'b11?????001001?????1?????????????,
                           TAimiatoo = 32'b11?????001001?????1?????????????,
                           CN = 32'b11?????001001?????1?????????????,
                           C = 32'b11?????001001?????1?????????????,
                           S = 32'b11?????001001?????1?????????????,
                           Si = 32'b11?????001001?????1?????????????,
                           Sami = 32'b11?????001001?????1?????????????,
                           Siami = 32'b11?????001001?????1?????????????,
                           Rs = 32'b11?????001001?????1?????????????,
                           Swc = 32'b11?????001001?????1?????????????,
                           Siwc = 32'b11?????001001?????1?????????????,
                           Swcami = 32'b11?????001001?????1?????????????,
                           Siwcami = 32'b11?????001001?????1?????????????,
                           Rswc = 32'b11?????001001?????1?????????????,
                           Tsami = 32'b11?????001001?????1?????????????,
                           Tsiami = 32'b11?????001001?????1?????????????,
                           Tsmiatoo = 32'b11?????001001?????1?????????????,
                           Tsimiatoo = 32'b11?????001001?????1?????????????,
                           BA = 32'b11?????001001?????1?????????????,
                           BA = 32'b11?????001001?????1?????????????,
                           BAamti = 32'b11?????001001?????1?????????????,
                           BAamti = 32'b11?????001001?????1?????????????,
                           BAwc = 32'b11?????001001?????1?????????????,
                           BAwc = 32'b11?????001001?????1?????????????,
                           BAwcami = 32'b11?????001001?????1?????????????,
                           BAwcami = 32'b11?????001001?????1?????????????,
                           BX = 32'b11?????001001?????1?????????????,
                           BX = 32'b11?????001001?????1?????????????,
                           BXamti = 32'b11?????001001?????1?????????????,
                           BXamti = 32'b11?????001001?????1?????????????,
                           BXwc = 32'b11?????001001?????1?????????????,
                           BXwc = 32'b11?????001001?????1?????????????,
                           BXwcami = 32'b11?????001001?????1?????????????,
                           BXwcami = 32'b11?????001001?????1?????????????,
                           BO = 32'b11?????001001?????1?????????????,
                           BO = 32'b11?????001001?????1?????????????,
                           BOamti = 32'b11?????001001?????1?????????????,
                           BOamti = 32'b11?????001001?????1?????????????,
                           BOwc = 32'b11?????001001?????1?????????????,
                           BOwc = 32'b11?????001001?????1?????????????,
                           BOwcami = 32'b11?????001001?????1?????????????,
                           BOwcami = 32'b11?????001001?????1?????????????,
                           Sll = 32'b11?????001001?????1?????????????,
                           Srl = 32'b11?????001001?????1?????????????,
                           Sra = 32'b11?????001001?????1?????????????,
                           Slli = 32'b11?????001001?????1?????????????,
                           Srli = 32'b11?????001001?????1?????????????,
                           Srai = 32'b11?????001001?????1?????????????,
                           JaL = 32'b11?????001001?????1?????????????,
                           JaLr = 32'b11?????001001?????1?????????????,
                           RfT = 32'b11?????001001?????1?????????????,
                           CaL = 32'b11?????001001?????1?????????????,
                           BN = 32'b11?????001001?????1?????????????,
                           BA = 32'b11?????001001?????1?????????????,
                           BTA = 32'b11?????001001?????1?????????????,
                           BAL = 32'b11?????001001?????1?????????????,
                           Bie = 32'b11?????001001?????1?????????????,
                           Bine = 32'b11?????001001?????1?????????????,
                           Bigtoe = 32'b11?????001001?????1?????????????,
                           Biltoe = 32'b11?????001001?????1?????????????,
                           Bigtoe( = 32'b11?????001001?????1?????????????,
                           Biltoe( = 32'b11?????001001?????1?????????????,
                           Bie( = 32'b11?????001001?????1?????????????,
                           Bine( = 32'b11?????001001?????1?????????????,
                           BoG = 32'b11?????001001?????1?????????????,
                           BoLoE = 32'b11?????001001?????1?????????????,
                           BoL = 32'b11?????001001?????1?????????????,
                           BoGU = 32'b11?????001001?????1?????????????,
                           BoCS(tU = 32'b11?????001001?????1?????????????,
                           BoP = 32'b11?????001001?????1?????????????,
                           BoN = 32'b11?????001001?????1?????????????,
                           BoOC = 32'b11?????001001?????1?????????????,
                           BoOS = 32'b11?????001001?????1?????????????,
                           Bo = 32'b11?????001001?????1?????????????,
                           C = 32'b11?????001001?????1?????????????,
                           CC = 32'b11?????001001?????1?????????????,
                           Sh2b = 32'b11?????001001?????1?????????????,
                           S( = 32'b11?????001001?????1?????????????,
                           Si( = 32'b11?????001001?????1?????????????,
                           R( = 32'b11?????001001?????1?????????????,
                           Ri( = 32'b11?????001001?????1?????????????,
                           trfc = 32'b11?????001001?????1?????????????,
                           tcfr = 32'b11?????001001?????1?????????????,
                           n = 32'b11?????001001?????1?????????????,
                           = 32'b11?????001001?????1?????????????,
                           RY = 32'b11?????001001?????1?????????????,
                           RP = 32'b11?????001001?????1?????????????,
                           Rw = 32'b11?????001001?????1?????????????,
                           Rt = 32'b11?????001001?????1?????????????,
                           Ra = 32'b11?????001001?????1?????????????,
                           WfrtY = 32'b11?????001001?????1?????????????,
                           WfitY = 32'b11?????001001?????1?????????????,
                           Wfrtp = 32'b11?????001001?????1?????????????,
                           Wfitp = 32'b11?????001001?????1?????????????,
                           Wfrtw = 32'b11?????001001?????1?????????????,
                           Wfitw = 32'b11?????001001?????1?????????????,
                           Wfrtt = 32'b11?????001001?????1?????????????,
                           Wfitt = 32'b11?????001001?????1?????????????,
                           wr,ra = 32'b11?????001001?????1?????????????,
                           Si = 32'b11?????001001?????1?????????????,
                           N = 32'b11?????001001?????1?????????????,
                           CO = 32'b11?????001001?????1?????????????,
                           CO = 32'b11?????001001?????1?????????????,
                           TA = 32'b11?????001001?????1?????????????,
                           TN = 32'b11?????001001?????1?????????????,
                           ToNE = 32'b11?????001001?????1?????????????,
                           ToE = 32'b11?????001001?????1?????????????,
                           ToG = 32'b11?????001001?????1?????????????,
                           ToLoE = 32'b11?????001001?????1?????????????,
                           ToGoE = 32'b11?????001001?????1?????????????,
                           ToL = 32'b11?????001001?????1?????????????,
                           ToGU = 32'b11?????001001?????1?????????????,
                           ToLoEU = 32'b11?????001001?????1?????????????,
                           ToCC(toEU = 32'b11?????001001?????1?????????????,
                           ToCS(TU = 32'b11?????001001?????1?????????????,
                           ToP = 32'b11?????001001?????1?????????????,
                           ToN = 32'b11?????001001?????1?????????????,
                           ToOC = 32'b11?????001001?????1?????????????,
                           ToOS = 32'b11?????001001?????1?????????????,
                           " = 32'b11?????001001?????1?????????????,
                           I = 32'b11?????001001?????1?????????????,
                           "I = 32'b11?????001001?????1?????????????,
                           = 32'b11?????001001?????1?????????????,


                            } opcode;
    `endif
endpackage